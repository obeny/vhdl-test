../../../src/bidir.vhd