../../../src/counter_gen.vhd