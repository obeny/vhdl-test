../../../src/and_gate.vhd