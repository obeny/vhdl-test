../../../src/xor_gate.vhd