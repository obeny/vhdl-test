../../../src/ff_d.vhd