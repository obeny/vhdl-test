../../../src/mux.vhd