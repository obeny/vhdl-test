../../../src/hiz_out.vhd